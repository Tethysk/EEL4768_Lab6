`include "muxes_a.v"
`include "muxes_b.v"
`include "muxes_c.v"

module mux21_tb;
reg wD0, wD1, wS;